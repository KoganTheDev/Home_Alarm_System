--------------------- Title ------------------------
-- Project Name: HA_System
-- File Name: Display_data.vhd
-- Author: Roni Shifrin
-- Ver: 0
-- Created Date: 23/11/25
----------------------------------------------------
