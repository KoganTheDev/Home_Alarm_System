--------------------- Title ------------------------
-- Project Name: HA_System
-- File Name: Code_register_TB.vhd
-- Author: Yuval Kogan
-- Ver: 0
-- Created Date: 23/11/25
----------------------------------------------------
